module main

const version = '0.0.0'
