module cmd

import cli

// https://github.com/opencontainers/runtime-spec/blob/master/runtime.md#create

fn create(command cli.Command) ? {
	println('Not implemented')
}
