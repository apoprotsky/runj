module cmd

import cli

fn start(cmd cli.Command) ? {
	println('Not implemented')
}
