module cmd

import cli

fn kill(cmd cli.Command) ? {
	println('Not implemented')
}
