module spec

pub const config = 'config.json'
