module cmd

import cli

fn state(cmd cli.Command) ? {
	println('Not implemented')
}
