module cmd

import cli

fn delete(cmd cli.Command) ? {
	println('Not implemented')
}
