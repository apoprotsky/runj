module state

const dir = '/var/db/runj/containers'
