module cmd

import cli

fn spec_command(command cli.Command) ? {
	println('Not implemented')
}
